// ysyx_22050710
module ysyx_22050710_clint (
  
);

  

endmodule
