// ysyx_22050710 Execute Unit csr
// ysyx_22050710
module ysyx_22050710_exu_csr (
  input [11:0] i_csraddr,
  input [4:0] i_rs1_or_zimm,
);

  

endmodule
