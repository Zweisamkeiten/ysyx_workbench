module prior_encode83(x, en, y);

endmodule
