// ysyx_22050710

module ysyx_22050710_if (
  input i_pc,
  output o_inst
);

  

endmodule
